

module add(input [7:0]DOut2,input [7:0]DOut1,output [7:0]ADDOut);


assign ADDOut = DOut2 + DOut1;    


endmodule
