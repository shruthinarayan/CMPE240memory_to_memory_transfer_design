


module sub(input [7:0]DOut2,input [7:0]DOut1,output [7:0]SUBOut);


assign SUBOut = DOut2 - DOut1;    


endmodule